module gpioTest(clock, out);

	input clock;
	output out;

	assign out = clock;

endmodule // gpioTest